module add_32(a,b,p);
  input [0:31] a,b;
  output [0:32] p;
  wire [0:31] s,c;
  assign p[0:31]=s[0:31];
  assign p[32]=c[31];
  add(a[0],b[0],0,c[0],s[0]);
  add(a[1],b[1],c[0],c[1],s[1]);
  add(a[2],b[2],c[1],c[2],s[2]);
  add(a[3],b[3],c[2],c[3],s[3]);
  add(a[4],b[4],c[3],c[4],s[4]);
  add(a[5],b[5],c[4],c[5],s[5]);
  add(a[6],b[6],c[5],c[6],s[6]);
  add(a[7],b[7],c[6],c[7],s[7]);
  add(a[8],b[8],c[7],c[8],s[8]);
  add(a[9],b[9],c[8],c[9],s[9]);
  add(a[10],b[10],c[9],c[10],s[10]);
  add(a[11],b[11],c[10],c[11],s[11]);
  add(a[12],b[12],c[11],c[12],s[12]);
  add(a[13],b[13],c[12],c[13],s[13]);
  add(a[14],b[14],c[13],c[14],s[14]);
  add(a[15],b[15],c[14],c[15],s[15]);
  add(a[16],b[16],c[15],c[16],s[16]);
  add(a[17],b[17],c[16],c[17],s[17]);
  add(a[18],b[18],c[17],c[18],s[18]);
  add(a[19],b[19],c[18],c[19],s[19]);
  add(a[20],b[20],c[19],c[20],s[20]);
  add(a[21],b[21],c[20],c[21],s[21]);
  add(a[22],b[22],c[21],c[22],s[22]);
  add(a[23],b[23],c[22],c[23],s[23]);
  add(a[24],b[24],c[23],c[24],s[24]);
  add(a[25],b[25],c[24],c[25],s[25]);
  add(a[26],b[26],c[25],c[26],s[26]);
  add(a[27],b[27],c[26],c[27],s[27]);
  add(a[28],b[28],c[27],c[28],s[28]);
  add(a[29],b[29],c[28],c[29],s[29]);
  add(a[30],b[30],c[29],c[30],s[30]);
  add(a[31],b[31],c[30],c[31],s[31]);
endmodule