module	mul5(f,m,p);
input	[4:0]	f,m;
output	[9:0]	p;
wire	[19:0]	s,c;
assign	p[0]=f[0]&m[0];
assign	{c[0],s[0]}=(f[1]&m[0])+(f[0]&m[1]);
assign	p[1]=s[0];
assign	{c[1],s[1]}=(f[2]&m[0])+(f[1]&m[1])+c[0];
assign	{c[2],s[2]}=(f[0]&m[2])+s[1];
assign	p[2]=s[2];
assign	{c[3],s[3]}=(f[3]&m[0])+(f[2]&m[1])+c[1];
assign	{c[4],s[4]}=(f[1]&m[2])+s[3]+c[2];
assign	{c[5],s[5]}=(f[0]&m[3])+s[4];
assign	p[3]=s[5];
assign	{c[6],s[6]}=(f[4]&m[0])+(f[3]&m[1])+c[3];
assign	{c[7],s[7]}=(f[2]&m[2])+s[6]+c[4];
assign	{c[8],s[8]}=(f[1]&m[3])+s[7]+c[5];
assign	{c[9],s[9]}=(f[0]&m[4])+s[8];
assign	p[4]=s[9];
assign	{c[10],s[10]}=(f[4]&m[1])+(f[3]&m[2])+c[6];
assign	{c[11],s[11]}=(f[2]&m[3])+s[10]+c[7];
assign	{c[12],s[12]}=(f[1]&m[4])+s[11]+c[8];
assign	{c[13],s[13]}=s[12]+c[9];
assign	p[5]=s[13];
assign	{c[14],s[14]}=(f[4]&m[2])+(f[3]&m[3])+c[10];
assign	{c[15],s[15]}=(f[2]&m[4])+s[14]+c[11];
assign	{c[16],s[16]}=s[15]+c[12]+c[13];
assign	p[6]=s[16];
assign	{c[17],s[17]}=(f[4]&m[3])+(f[3]&m[4])+c[14];
assign	{c[18],s[18]}=s[17]+c[15]+c[16];
assign	p[7]=s[18];
assign	{c[19],s[19]}=(f[4]&m[4])+c[17]+c[18];
assign	p[8]=s[19];
assign	p[9]=c[19];
endmodule