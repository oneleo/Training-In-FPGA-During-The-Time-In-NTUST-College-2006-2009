module print_7(z,p);
  input [3:0] z;
  output [6:0] p;
  assign p[0]=~z[3]&~z[2]&~z[1]&~z[0] | ~z[3]&~z[2]&z[1]&~z[0] | ~z[3]&~z[2]&z[1]&z[0] | ~z[3]&z[2]&~z[1]&z[0] | ~z[3]&z[2]&z[1]&~z[0] | ~z[3]&z[2]&z[1]&z[0] | z[3]&~z[2]&~z[1]&~z[0] | z[3]&~z[2]&~z[1]&z[0] | z[3]&~z[2]&z[1]&~z[0] | z[3]&z[2]&~z[1]&~z[0] | z[3]&z[2]&z[1]&~z[0] | z[3]&z[2]&z[1]&z[0];
  assign p[1]=~z[3]&~z[2]&~z[1]&~z[0] | ~z[3]&~z[2]&~z[1]&z[0] | ~z[3]&~z[2]&z[1]&~z[0] | ~z[3]&~z[2]&z[1]&z[0] | ~z[3]&z[2]&~z[1]&~z[0] | ~z[3]&z[2]&z[1]&z[0] | z[3]&~z[2]&~z[1]&~z[0] | z[3]&~z[2]&~z[1]&z[0] | z[3]&~z[2]&z[1]&~z[0] | z[3]&z[2]&~z[1]&z[0];
  assign p[2]=~z[3]&~z[2]&~z[1]&~z[0] | ~z[3]&~z[2]&~z[1]&z[0] | ~z[3]&~z[2]&z[1]&z[0] | ~z[3]&z[2]&~z[1]&~z[0] | ~z[3]&z[2]&~z[1]&z[0] | ~z[3]&z[2]&z[1]&~z[0] | ~z[3]&z[2]&z[1]&z[0] | z[3]&~z[2]&~z[1]&~z[0] | z[3]&~z[2]&~z[1]&z[0] | z[3]&~z[2]&z[1]&z[0] | z[3]&z[2]&~z[1]&z[0]; 
  assign p[3]=~z[3]&~z[2]&~z[1]&~z[0] | ~z[3]&~z[2]&z[1]&~z[0] | ~z[3]&~z[2]&z[1]&z[0] | ~z[3]&z[2]&~z[1]&z[0] | ~z[3]&z[2]&z[1]&~z[0] | z[3]&~z[2]&~z[1]&~z[0] | z[3]&~z[2]&~z[1]&z[0] | z[3]&~z[2]&z[1]&~z[0] | z[3]&~z[2]&z[1]&z[0] | z[3]&z[2]&~z[1]&~z[0] | z[3]&z[2]&~z[1]&z[0] | z[3]&z[2]&z[1]&~z[0];
  assign p[4]=~z[3]&~z[2]&~z[1]&~z[0] | ~z[3]&~z[2]&z[1]&~z[0] | ~z[3]&z[2]&z[1]&~z[0] | z[3]&~z[2]&~z[1]&~z[0] | z[3]&~z[2]&z[1]&~z[0] | z[3]&~z[2]&z[1]&z[0] | z[3]&z[2]&~z[1]&~z[0] | z[3]&z[2]&~z[1]&z[0] | z[3]&z[2]&z[1]&~z[0] | z[3]&z[2]&z[1]&z[0];
  assign p[5]=~z[3]&~z[2]&~z[1]&~z[0] | ~z[3]&z[2]&~z[1]&~z[0] | ~z[3]&z[2]&~z[1]&z[0] | ~z[3]&z[2]&z[1]&~z[0] | z[3]&~z[2]&~z[1]&~z[0] | z[3]&~z[2]&~z[1]&z[0] | z[3]&~z[2]&z[1]&~z[0] | z[3]&~z[2]&z[1]&z[0] | z[3]&z[2]&~z[1]&~z[0] | z[3]&z[2]&z[1]&~z[0] | z[3]&z[2]&z[1]&z[0];
  assign p[6]=~z[3]&~z[2]&z[1]&~z[0] | ~z[3]&~z[2]&z[1]&z[0] | ~z[3]&z[2]&~z[1]&~z[0] | ~z[3]&z[2]&~z[1]&z[0] | ~z[3]&z[2]&z[1]&~z[0] | z[3]&~z[2]&~z[1]&~z[0] | z[3]&~z[2]&~z[1]&z[0] | z[3]&~z[2]&z[1]&~z[0] | z[3]&~z[2]&z[1]&z[0] | z[3]&z[2]&~z[1]&z[0] | z[3]&z[2]&z[1]&~z[0] | z[3]&z[2]&z[1]&z[0];
endmodule