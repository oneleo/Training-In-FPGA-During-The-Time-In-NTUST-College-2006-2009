/*module print_7(z,a,b,c,d,e,f,g);
  input [3:0] z;
  output a,b,c,d,e,f,g;
  assign a=~z[3]&~z[2]&~z[1]&~z[0] | ~z[3]&~z[2]&z[1]&~z[0] | ~z[3]&~z[2]&z[1]&z[0] | ~z[3]&z[2]&~z[1]&z[0] | ~z[3]&z[2]&z[1]&~z[0] | ~z[3]&z[2]&z[1]&z[0] | z[3]&~z[2]&~z[1]&~z[0] | z[3]&~z[2]&~z[1]&z[0] | z[3]&~z[2]&z[1]&~z[0] | z[3]&z[2]&~z[1]&~z[0] | z[3]&z[2]&z[1]&~z[0] | z[3]&z[2]&z[1]&z[0];
  assign b=~z[3]&~z[2]&~z[1]&~z[0] | ~z[3]&~z[2]&~z[1]&z[0] | ~z[3]&~z[2]&z[1]&~z[0] | ~z[3]&~z[2]&z[1]&z[0] | ~z[3]&z[2]&~z[1]&~z[0] | ~z[3]&z[2]&z[1]&z[0] | z[3]&~z[2]&~z[1]&~z[0] | z[3]&~z[2]&~z[1]&z[0] | z[3]&~z[2]&z[1]&~z[0] | z[3]&z[2]&~z[1]&z[0];
  assign c=~z[3]&~z[2]&~z[1]&~z[0] | ~z[3]&~z[2]&~z[1]&z[0] | ~z[3]&~z[2]&z[1]&z[0] | ~z[3]&z[2]&~z[1]&~z[0] | ~z[3]&z[2]&~z[1]&z[0] | ~z[3]&z[2]&z[1]&~z[0] | ~z[3]&z[2]&z[1]&z[0] | z[3]&~z[2]&~z[1]&~z[0] | z[3]&~z[2]&~z[1]&z[0] | z[3]&~z[2]&z[1]&z[0] | z[3]&z[2]&~z[1]&z[0]; 
  assign d=~z[3]&~z[2]&~z[1]&~z[0] | ~z[3]&~z[2]&z[1]&~z[0] | ~z[3]&~z[2]&z[1]&z[0] | ~z[3]&z[2]&~z[1]&z[0] | ~z[3]&z[2]&z[1]&~z[0] | z[3]&~z[2]&~z[1]&~z[0] | z[3]&~z[2]&~z[1]&z[0] | z[3]&~z[2]&z[1]&~z[0] | z[3]&~z[2]&z[1]&z[0] | z[3]&z[2]&~z[1]&~z[0] | z[3]&z[2]&~z[1]&z[0] | z[3]&z[2]&z[1]&~z[0];
  assign e=~z[3]&~z[2]&~z[1]&~z[0] | ~z[3]&~z[2]&z[1]&~z[0] | ~z[3]&z[2]&z[1]&~z[0] | z[3]&~z[2]&~z[1]&~z[0] | z[3]&~z[2]&z[1]&~z[0] | z[3]&~z[2]&z[1]&z[0] | z[3]&z[2]&~z[1]&~z[0] | z[3]&z[2]&~z[1]&z[0] | z[3]&z[2]&z[1]&~z[0] | z[3]&z[2]&z[1]&z[0];
  assign f=~z[3]&~z[2]&~z[1]&~z[0] | ~z[3]&z[2]&~z[1]&~z[0] | ~z[3]&z[2]&~z[1]&z[0] | ~z[3]&z[2]&z[1]&~z[0] | z[3]&~z[2]&~z[1]&~z[0] | z[3]&~z[2]&~z[1]&z[0] | z[3]&~z[2]&z[1]&~z[0] | z[3]&~z[2]&z[1]&z[0] | z[3]&z[2]&~z[1]&~z[0] | z[3]&z[2]&z[1]&~z[0] | z[3]&z[2]&z[1]&z[0];
  assign g=~z[3]&~z[2]&z[1]&~z[0] | ~z[3]&~z[2]&z[1]&z[0] | ~z[3]&z[2]&~z[1]&~z[0] | ~z[3]&z[2]&~z[1]&z[0] | ~z[3]&z[2]&z[1]&~z[0] | z[3]&~z[2]&~z[1]&~z[0] | z[3]&~z[2]&~z[1]&z[0] | z[3]&~z[2]&z[1]&~z[0] | z[3]&~z[2]&z[1]&z[0] | z[3]&z[2]&~z[1]&z[0] | z[3]&z[2]&z[1]&~z[0] | z[3]&z[2]&z[1]&z[0];
endmodule*/
module print_7(z,a,b,c,d,e,f,g);
  input [3:0] z;
  output a,b,c,d,e,f,g;
  assign a=(z==0)|(z==2)|(z==3)|(z==5)|(z==6)|(z==7)|(z==8)|(z==9)|(z==10)|(z==12)|(z==14)|(z==15);
  assign b=(z==0)|(z==1)|(z==2)|(z==3)|(z==4)|(z==7)|(z==8)|(z==9)|(z==10)|(z==13);
  assign c=(z==0)|(z==1)|(z==3)|(z==4)|(z==5)|(z==6)|(z==7)|(z==8)|(z==9)|(z==11)|(z==13);
  assign d=(z==0)|(z==2)|(z==3)|(z==5)|(z==6)|(z==8)|(z==9)|(z==10)|(z==11)|(z==12)|(z==13)|(z==14);
  assign e=(z==0)|(z==2)|(z==6)|(z==8)|(z==10)|(z==11)|(z==12)|(z==13)|(z==14)|(z==15);
  assign f=(z==0)|(z==4)|(z==5)|(z==6)|(z==8)|(z==9)|(z==10)|(z==11)|(z==12)|(z==14)|(z==15);
  assign g=(z==2)|(z==3)|(z==4)|(z==5)|(z==6)|(z==8)|(z==9)|(z==10)|(z==11)|(z==13)|(z==14)|(z==15);
endmodule